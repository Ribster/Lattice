LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY lattice;
USE work.constants.all;

package functions is

end functions;

package body functions is

end functions;