LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY lattice;
USE work.constants.all;

package functions is
	-- function prototypes
	function to_std_logic(arg : boolean) return std_logic; 
	function to_boolean(arg: std_logic) return boolean;
	function hstr(slv: std_logic_vector) return string;
end functions;

package body functions is
	--
	-- convert a boolean to a std_logic
	--
	function to_std_logic(arg : boolean) return std_logic is 
	begin 
		if arg then 
		  return '1'; 
		else 
		  return '0'; 
		end if; 
	end function to_std_logic;

	--
	-- convert a std_logic to a boolean
	--
	function to_boolean(arg : std_logic) return boolean is
	begin
		if arg = '1' then
		  return true;
		else
		  return false;
		end if;
	end function to_boolean;

	-- 
	-- useful hex converter for simulation reporting only
	--
	function hstr(slv: std_logic_vector) return string is
		variable hexlen: integer;
		variable longslv : std_logic_vector(67 downto 0) := (others => '0');
		variable hex : string(1 to 20);
		variable fourbit : std_logic_vector(3 downto 0);
		begin
			hexlen := (slv'left+1)/4;
			
			if (slv'left+1) mod 4 /= 0 then
			 hexlen := hexlen + 1;
			end if;
			
			longslv(slv'left downto 0) := slv;
			
			for i in (hexlen -1) downto 0 loop
			 fourbit := longslv(((i*4)+3) downto (i*4));
				 case fourbit is
				   when "0000" => hex(hexlen -I) := '0';
				   when "0001" => hex(hexlen -I) := '1';
				   when "0010" => hex(hexlen -I) := '2';
				   when "0011" => hex(hexlen -I) := '3';
				   when "0100" => hex(hexlen -I) := '4';
				   when "0101" => hex(hexlen -I) := '5';
				   when "0110" => hex(hexlen -I) := '6';
				   when "0111" => hex(hexlen -I) := '7';
				   when "1000" => hex(hexlen -I) := '8';
				   when "1001" => hex(hexlen -I) := '9';
				   when "1010" => hex(hexlen -I) := 'A';
				   when "1011" => hex(hexlen -I) := 'B';
				   when "1100" => hex(hexlen -I) := 'C';
				   when "1101" => hex(hexlen -I) := 'D';
				   when "1110" => hex(hexlen -I) := 'E';
				   when "1111" => hex(hexlen -I) := 'F';
				   when "ZZZZ" => hex(hexlen -I) := 'z';
				   when "UUUU" => hex(hexlen -I) := 'u';
				   when "XXXX" => hex(hexlen -I) := 'x';
				   when others => hex(hexlen -I) := '?';
				 end case;
			end loop;
		return hex(1 to hexlen);
	end hstr;

end functions;